CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
75 C:\Users\Adrianne\AppData\Local\Temp\Rar$EXa0.190\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
30
13 Logic Switch~
5 41 322 0 10 11
0 16 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3409 0 0
2
42879.3 0
0
13 Logic Switch~
5 40 283 0 10 11
0 18 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3951 0 0
2
42879.3 1
0
13 Logic Switch~
5 38 242 0 10 11
0 20 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8885 0 0
2
42879.3 2
0
13 Logic Switch~
5 40 202 0 10 11
0 19 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3780 0 0
2
42879.3 3
0
13 Logic Switch~
5 35 164 0 10 11
0 23 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9265 0 0
2
42879.3 4
0
13 Logic Switch~
5 37 129 0 1 11
0 22
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9442 0 0
2
42879.3 5
0
13 Logic Switch~
5 35 92 0 10 11
0 26 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9424 0 0
2
42879.3 6
0
13 Logic Switch~
5 36 50 0 10 11
0 25 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9968 0 0
2
42879.3 7
0
2 +V
167 299 670 0 1 3
0 3
0
0 0 54256 0
3 10V
-11 -22 10 -14
3 V11
-11 -32 10 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9281 0 0
2
5.89801e-315 0
0
2 +V
167 252 670 0 1 3
0 4
0
0 0 54256 0
3 10V
-11 -22 10 -14
3 V10
-11 -32 10 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8464 0 0
2
5.89801e-315 0
0
2 +V
167 196 669 0 1 3
0 5
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V9
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7168 0 0
2
5.89801e-315 0
0
14 Logic Display~
6 589 478 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3171 0 0
2
42879.3 8
0
14 Logic Display~
6 654 311 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4139 0 0
2
42879.3 9
0
14 Logic Display~
6 596 150 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6435 0 0
2
42879.3 10
0
5 4001~
219 599 329 0 3 22
0 2 7 6
0
0 0 624 0
4 4001
-14 -24 14 -16
3 U8A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 7 0
1 U
5283 0 0
2
42879.3 11
0
8 4-In OR~
219 488 497 0 5 22
0 11 10 9 8 7
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U7A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 6 0
1 U
6874 0 0
2
42879.3 12
0
5 4049~
219 135 588 0 2 22
0 16 17
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U4E
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 4 0
1 U
5305 0 0
2
42879.3 13
0
5 4049~
219 243 507 0 2 22
0 20 21
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U4D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 4 0
1 U
34 0 0
2
42879.3 14
0
5 4049~
219 417 592 0 2 22
0 12 8
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U4C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 4 0
1 U
969 0 0
2
42879.3 15
0
5 4068~
219 368 592 0 9 19
0 13 14 15 17 18 5 4 3 12
0
0 0 624 0
4 4068
-7 -24 21 -16
2 U6
-8 -44 6 -36
0
15 DVDD=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 2 3 4 5 9 10 11 12 13
2 3 4 5 9 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
8402 0 0
2
42879.3 16
0
5 4082~
219 364 503 0 5 22
0 13 14 21 19 9
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U2B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 2 0
1 U
3751 0 0
2
42879.3 17
0
5 4049~
219 244 441 0 2 22
0 23 24
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U4B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 4 0
1 U
4292 0 0
2
42879.3 18
0
5 4073~
219 361 442 0 4 22
0 13 24 22 10
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 5 0
1 U
6118 0 0
2
42879.3 19
0
5 4049~
219 240 372 0 2 22
0 26 27
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U4A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 4 0
1 U
34 0 0
2
42879.3 20
0
5 4081~
219 358 381 0 3 22
0 27 25 11
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 3 0
1 U
6357 0 0
2
42879.3 21
0
5 4082~
219 408 175 0 5 22
0 13 14 15 28 2
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U2A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 2 0
1 U
319 0 0
2
42879.3 22
0
10 2-In XNOR~
219 227 299 0 3 22
0 18 16 28
0
0 0 624 0
4 4077
-7 -24 21 -16
3 U1D
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 1 0
1 U
3976 0 0
2
42879.3 23
0
10 2-In XNOR~
219 229 216 0 3 22
0 19 20 15
0
0 0 624 0
4 4077
-7 -24 21 -16
3 U1C
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 1 0
1 U
7634 0 0
2
42879.3 24
0
10 2-In XNOR~
219 226 139 0 3 22
0 22 23 14
0
0 0 624 0
4 4077
-7 -24 21 -16
3 U1B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 1 0
1 U
523 0 0
2
42879.3 25
0
10 2-In XNOR~
219 225 74 0 3 22
0 25 26 13
0
0 0 624 0
4 4077
-7 -24 21 -16
3 U1A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
6748 0 0
2
42879.3 26
0
43
1 0 2 0 0 8192 0 15 0 0 2 3
586 320
560 320
560 175
5 1 2 0 0 4224 0 26 14 0 0 3
429 175
596 175
596 168
1 8 3 0 0 8320 0 9 20 0 0 4
299 679
314 679
314 624
344 624
1 7 4 0 0 12416 0 10 20 0 0 4
252 679
269 679
269 615
344 615
1 6 5 0 0 12416 0 11 20 0 0 4
196 678
222 678
222 606
344 606
3 1 6 0 0 4224 0 15 13 0 0 2
638 329
654 329
0 1 7 0 0 4096 0 0 12 8 0 2
560 496
589 496
5 2 7 0 0 8336 0 16 15 0 0 4
521 497
560 497
560 338
586 338
2 4 8 0 0 12416 0 19 16 0 0 5
438 592
438 594
437 594
437 511
471 511
5 3 9 0 0 4224 0 21 16 0 0 3
385 503
471 503
471 502
4 2 10 0 0 4224 0 23 16 0 0 4
382 442
437 442
437 493
471 493
3 1 11 0 0 8320 0 25 16 0 0 4
379 381
454 381
454 484
471 484
9 1 12 0 0 4224 0 20 19 0 0 4
395 592
403 592
403 592
402 592
1 0 13 0 0 8320 0 20 0 0 35 3
344 561
332 561
332 74
2 0 14 0 0 8320 0 20 0 0 34 3
344 570
320 570
320 139
3 0 15 0 0 8320 0 20 0 0 33 3
344 579
309 579
309 216
1 0 16 0 0 8320 0 17 0 0 36 3
120 588
96 588
96 308
2 4 17 0 0 4224 0 17 20 0 0 2
156 588
344 588
5 0 18 0 0 8320 0 20 0 0 37 3
344 597
114 597
114 290
4 0 19 0 0 8320 0 21 0 0 39 3
340 517
129 517
129 207
1 0 20 0 0 8320 0 18 0 0 38 3
228 507
145 507
145 225
2 0 14 0 0 0 0 21 0 0 34 3
340 499
297 499
297 139
1 0 13 0 0 0 0 21 0 0 35 3
340 490
287 490
287 74
2 3 21 0 0 8320 0 18 21 0 0 3
264 507
264 508
340 508
3 0 22 0 0 8320 0 23 0 0 41 3
337 451
158 451
158 139
1 0 23 0 0 8320 0 22 0 0 40 3
229 441
172 441
172 148
2 2 24 0 0 8320 0 22 23 0 0 3
265 441
265 442
337 442
1 0 13 0 0 0 0 23 0 0 35 3
337 433
273 433
273 74
2 0 25 0 0 8320 0 25 0 0 43 3
334 390
184 390
184 65
1 0 26 0 0 8320 0 24 0 0 42 3
225 372
196 372
196 83
2 1 27 0 0 12416 0 24 25 0 0 4
261 372
259 372
259 372
334 372
3 4 28 0 0 8320 0 27 26 0 0 4
266 299
363 299
363 189
384 189
3 3 15 0 0 0 0 28 26 0 0 4
268 216
344 216
344 180
384 180
3 2 14 0 0 0 0 29 26 0 0 4
265 139
343 139
343 171
384 171
3 1 13 0 0 0 0 30 26 0 0 4
264 74
361 74
361 162
384 162
1 2 16 0 0 0 0 1 27 0 0 4
53 322
79 322
79 308
211 308
1 1 18 0 0 0 0 2 27 0 0 5
52 283
52 282
77 282
77 290
211 290
1 2 20 0 0 0 0 3 28 0 0 5
50 242
50 241
76 241
76 225
213 225
1 1 19 0 0 0 0 4 28 0 0 5
52 202
52 199
76 199
76 207
213 207
1 2 23 0 0 0 0 5 29 0 0 4
47 164
75 164
75 148
210 148
1 1 22 0 0 0 0 6 29 0 0 6
49 129
49 124
76 124
76 139
210 139
210 130
1 2 26 0 0 0 0 7 30 0 0 4
47 92
76 92
76 83
209 83
1 1 25 0 0 0 0 8 30 0 0 4
48 50
76 50
76 65
209 65
11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
591 470 652 494
601 478 641 494
5 A > B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
660 306 721 330
670 314 710 330
5 A < B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
598 154 659 178
608 162 648 178
5 A = B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
-7 306 30 330
3 314 19 330
2 B0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
-8 266 29 290
2 274 18 290
2 A0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
-8 225 29 249
2 233 18 249
2 B1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
-8 188 29 212
2 196 18 212
2 A1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
-9 149 28 173
1 157 17 173
2 B2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
-9 112 28 136
1 120 17 136
2 A2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
-6 77 31 101
4 85 20 101
2 B3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
-7 31 30 55
3 39 19 55
2 A3
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
